module hazard(
	input wire memread,
	input wire [4:0] rt_now,
	input wire [4:0] rs_now,
	input wire [4:0] rt_pre,
	input wire [4:0] rs_pre,
	output reg stall

);

	// {{{ load use data hazard detection, signal stall

	/* If an operation in stage 4 (MEM) loads from memory (e.g. lw)
	 * and the operation in stage 3 (EX) depends on this value,
	 * a stall must be performed.  The memory read cannot 
	 * be forwarded because memory access is too slow.  It can
	 * be forwarded from stage 5 (WB) after a stall.
	 *
	 *   lw $1, 16($10)  ; I-type, rt_s3 = $1, memread_s3 = 1
	 *   sw $1, 32($12)  ; I-type, rt_s2 = $1, memread_s2 = 0
	 *
	 *   lw $1, 16($3)  ; I-type, rt_s3 = $1, memread_s3 = 1
	 *   sw $2, 32($1)  ; I-type, rt_s2 = $2, rs_s2 = $1, memread_s2 = 0
	 *
	 *   lw  $1, 16($3)  ; I-type, rt_s3 = $1, memread_s3 = 1
	 *   add $2, $1, $1  ; R-type, rs_s2 = $1, rt_s2 = $1, memread_s2 = 0
	 */
	
	always @(*) begin
		if (memread == 1'b1 && ((rt_now == rt_pre) || (rs_now == rt_pre)) ) begin
			stall <= 1'b1;  // perform a stall
		end else
			stall <= 1'b0;  // no stall
	end
	// }}}
endmodule
